*** Fund. de Projeto Analógico
** Caracterização NMOS e PMOS para 
** projeto gm/Id

*** Opcoes
** salvar as correntes para poder mostrar depois
.options savecurrents
.options filetype=ascii
.temp 25


** transistores
Mn vdd1 vg1 gnd gnd nmos l={2*lambda} w={20*lambda} ad={6*lambda*w} as={6*lambda*w} pd={12*lambda+2*w} ps={12*lambda+2*w}
Mp vdd2 vg2 gnd gnd pmos l={2*lambda} w={20*lambda} ad={6*lambda*w} as={6*lambda*w} pd={12*lambda+2*w} ps={12*lambda+2*w}

*** Parametros e Inclusoes
.include ../modelos_spice/130nm_bulk.pm
.param lambda=65n
.param w=20*lambda
.param vd=1.3
.param vg=0.3
.csparam vddsim={vd}

vdd vdd gnd dc vd
vgg vgg gnd dc vg

bdd1 vdd1 gnd v = v(vdd)
bdd2 vdd2 gnd v = '-v(vdd)'

bgg2 gnd vg2 v = v(vgg)
bgg1 vg1 gnd v = v(vgg)

*.dc vgg 0.7 1.5 0.01
*.dc vdd 0 5 10m
*.pz vg1 gnd vdd1 gnd pz
*.pz vg2 gnd vdd2 gnd pz
*.ac dec 100 1 1k

.end

.control
** Ajuste de opcoes
set color0=white
set color1=black
set units = degrees
set wr_singlescale
set wr_vecnames
set width = 4098
set filetype = ascii
*set appendwrite

** Parametros a serem salvos
save all @mn[id] @mn[ibs] @mn[gm] @mn[gds] @mn[gmbs] @mn[vdsat] @mn[vth]
				+@mn[cgs] @mn[cgd] @mn[cgb] @mn[cbd] @mn[cbs] 
        +@mn[cdd] @mn[cgg] @mn[css] @mn[cbb] @mn[capbd] @mn[capbs]
				+@mn[vgs] @mn[vds] @mn[vbs]
				+@mp[id] @mp[ibs] @mp[gm] @mp[gds] @mp[gmbs] @mp[vdsat] @mp[vth]
				+@mp[cgs] @mp[cgd] @mp[cgb] @mp[cbd] @mp[cbs] 
        +@mp[cdd] @mp[cgg] @mp[css] @mp[cbb] @mp[capbd] @mp[capbs]
				+@mp[vgs] @mp[vds] @mp[vbs]

*** Roda as simulacoes, calcula os parametros e salva em arquivo

* Cria as variaveis para fazer as simulacoes
let comp = 130n
let delta = 10n

* Loop para variar o comprimento de canal e 
while comp < 270n
	echo "Realizando simulação variando tensão na porta (Vgg) para L="$&comp"."
  * Modifica o comprimento dos transistores para o valor ajustado
	alter @mn[l] = comp 
  alter @mp[l] = comp
  * Realiza a simulacao CC variando a tensao de porta
	dc vgg 0 1.3 0.25m
  * Grava o comprimento para compor o nome do arquivo de saida
  let comp_ext = comp/1e-9
  * Incrementa o comprimento para a proxima simulacao
 	let comp = comp + delta

  * Tratamento de dados para os NMOS. A maioria eh soh exemplo.
  * Nao serao necessariamente usados.
  let mn.id			= @mn[id]
  let mn.ibs		= @mn[ibs]
  let mn.gm			= @mn[gm]
  let mn.gds		= @mn[gds]
  let mn.gmbs		= @mn[gmbs]
  let mn.vsat		= @mn[vdsat]
  let mn.vth    = @mn[vth]
  let mn.cgs		= @mn[cgs]
  let mn.cgd		= @mn[cgd]
  let mn.cgb		= @mn[cgb]
  let mn.cbd		= @mn[cbd]
  let mn.cbs		= @mn[cbs]
  let mn.cdd    = @mn[cdd] 
  let mn.cgg    = @mn[cgg] 
  let mn.css    = @mn[css] 
  let mn.cbb    = @mn[cbb] 
  let mn.capbd  = @mn[capbd] 
  let mn.capbs  = @mn[capbs]
  let mn.vgs		= @mn[vgs]
  let mn.vds		= @mn[vds]
  let mn.vbs		= @mn[vbs]
  let eff_n     = 'mn.gm/mn.id'
  let ov_n      = 'mn.vgs - mn.vth'
  let pi_2      = '2*3.14159'
  let ft_n      = '(1/pi_2)*(mn.gm/mn.cgg)'
  let av_n      = 'mn.gm/mn.gds'
  let id_w_n    = 'mn.id/@mn[w]'
  let ro_n      = '1/mn.gds'
  let eff_ft_n  = 'eff_n*ft_n'

  * Tratamento de dados para os PMOS
  let mp.id			= @mp[id]
  let mp.ibs		= @mp[ibs]
  let mp.gm			= @mp[gm]
  let mp.gds		= @mp[gds]
  let mp.gmbs		= @mp[gmbs]
  let mp.vsat		= @mp[vdsat]
  let mp.vth    = @mp[vth]
  let mp.cgs		= @mp[cgs]
  let mp.cgd		= @mp[cgd]
  let mp.cgb		= @mp[cgb]
  let mp.cbd		= @mp[cbd]
  let mp.cbs		= @mp[cbs]
  let mp.cdd    = @mp[cdd] 
  let mp.cgg    = @mp[cgg] 
  let mp.css    = @mp[css] 
  let mp.cbb    = @mp[cbb] 
  let mp.capbd  = @mp[capbd] 
  let mp.capbs  = @mp[capbs]
  let mp.vgs		= @mp[vgs]
  let mp.vds		= @mp[vds]
  let mp.vbs		= @mp[vbs]
  let eff_p     = 'mp.gm/mp.id'
  let ov_p      = 'mp.vgs - mp.vth'
  let ft_p      = '(1/pi_2)*(mp.gm/mp.cgg)'
  let av_p      = 'mp.gm/mp.gds'
  let id_w_p    = 'mp.id/@mp[w]'
  let ro_p      = '1/mp.gds'
  let eff_ft_p  = 'eff_p*ft_p'

  * Compoe o nome do arquivo para escrita. Extensao eh livre.
  set arquivo1	=	{'curvas_nmos_l_'}{$&comp_ext}{'n_vdd_'}{$&vddsim}{'.dat'}
  * Escreve os dados selecionados no arquivo
  wrdata $arquivo1	mn.id mn.gm mn.gds mn.gmbs mn.vsat mn.vth
                +mn.cgd mn.cgg mn.vgs mn.vds mn.vbs
                +eff_n ov_n ft_n av_n id_w_n ro_n eff_ft_n

  * Mesma coisa para os PMOS
  set arquivo2	=	{'curvas_pmos_l_'}{$&comp_ext}{'n_vdd_'}{$&vddsim}{'.dat'}
  wrdata $arquivo2	mp.id mp.gm mp.gds mp.gmbs mp.vsat mp.vth
                +mp.cgd mp.cgg mp.vgs mp.vds mp.vbs
                +eff_p ov_p ft_p av_p id_w_p ro_p eff_ft_p
end

plot dc1.eff_n dc2.eff_n dc3.eff_n dc4.eff_n dc5.eff_n dc6.eff_n dc7.eff_n dc8.eff_n dc9.eff_n dc10.eff_n dc11.eff_n dc12.eff_n dc13.eff_n dc14.eff_n

plot dc1.av_n vs dc1.eff_n dc2.av_n vs dc2.eff_n dc3.av_n vs dc3.eff_n dc4.av_n vs dc4.eff_n dc5.av_n vs dc5.eff_n dc6.av_n vs dc6.eff_n dc7.av_n vs dc7.eff_n dc8.av_n vs dc8.eff_n dc9.av_n vs dc9.eff_n dc10.av_n vs dc10.eff_n dc11.av_n vs dc11.eff_n dc12.av_n vs dc12.eff_n dc13.av_n vs dc13.eff_n dc14.av_n vs dc14.eff_n

plot dc1.ft_n vs dc1.eff_n dc2.ft_n vs dc2.eff_n dc3.ft_n vs dc3.eff_n dc4.ft_n vs dc4.eff_n dc5.ft_n vs dc5.eff_n dc6.ft_n vs dc6.eff_n dc7.ft_n vs dc7.eff_n dc8.ft_n vs dc8.eff_n dc9.ft_n vs dc9.eff_n dc10.ft_n vs dc10.eff_n dc11.ft_n vs dc11.eff_n dc12.ft_n vs dc12.eff_n dc13.ft_n vs dc13.eff_n dc14.ft_n vs dc14.eff_n

plot dc1.id_w_n vs dc1.eff_n ylog dc2.id_w_n vs dc2.eff_n dc3.id_w_n vs dc3.eff_n dc4.id_w_n vs dc4.eff_n dc5.id_w_n vs dc5.eff_n dc6.id_w_n vs dc6.eff_n dc7.id_w_n vs dc7.eff_n dc8.id_w_n vs dc8.eff_n dc9.id_w_n vs dc9.eff_n dc10.id_w_n vs dc10.eff_n dc11.id_w_n vs dc11.eff_n dc12.id_w_n vs dc12.eff_n dc13.id_w_n vs dc13.eff_n dc14.id_w_n vs dc14.eff_n

plot dc1.eff_ft_n vs dc1.eff_n dc2.eff_ft_n vs dc2.eff_n dc3.eff_ft_n vs dc3.eff_n dc4.eff_ft_n vs dc4.eff_n dc5.eff_ft_n vs dc5.eff_n dc6.eff_ft_n vs dc6.eff_n dc7.eff_ft_n vs dc7.eff_n dc8.eff_ft_n vs dc8.eff_n dc9.eff_ft_n vs dc9.eff_n dc10.eff_ft_n vs dc10.eff_n dc11.eff_ft_n vs dc11.eff_n dc12.eff_ft_n vs dc12.eff_n dc13.eff_ft_n vs dc13.eff_n dc14.eff_ft_n vs dc14.eff_n



plot dc1.eff_p dc2.eff_p dc3.eff_p dc4.eff_p dc5.eff_p dc6.eff_p dc7.eff_p dc8.eff_p dc9.eff_p dc10.eff_p dc11.eff_p dc12.eff_p dc13.eff_p dc14.eff_p

plot dc1.av_p vs dc1.eff_p dc2.av_p vs dc2.eff_p dc3.av_p vs dc3.eff_p dc4.av_p vs dc4.eff_p dc5.av_p vs dc5.eff_p dc6.av_p vs dc6.eff_p dc7.av_p vs dc7.eff_p dc8.av_p vs dc8.eff_p dc9.av_p vs dc9.eff_p dc10.av_p vs dc10.eff_p dc11.av_p vs dc11.eff_p dc12.av_p vs dc12.eff_p dc13.av_p vs dc13.eff_p dc14.av_p vs dc14.eff_p

plot dc1.ft_p vs dc1.eff_p dc2.ft_p vs dc2.eff_p dc3.ft_p vs dc3.eff_p dc4.ft_p vs dc4.eff_p dc5.ft_p vs dc5.eff_p dc6.ft_p vs dc6.eff_p dc7.ft_p vs dc7.eff_p dc8.ft_p vs dc8.eff_p dc9.ft_p vs dc9.eff_p dc10.ft_p vs dc10.eff_p dc11.ft_p vs dc11.eff_p dc12.ft_p vs dc12.eff_p dc13.ft_p vs dc13.eff_p dc14.ft_p vs dc14.eff_p

plot dc1.id_w_p vs dc1.eff_p ylog dc2.id_w_p vs dc2.eff_p dc3.id_w_p vs dc3.eff_p dc4.id_w_p vs dc4.eff_p dc5.id_w_p vs dc5.eff_p dc6.id_w_p vs dc6.eff_p dc7.id_w_p vs dc7.eff_p dc8.id_w_p vs dc8.eff_p dc9.id_w_p vs dc9.eff_p dc10.id_w_p vs dc10.eff_p dc11.id_w_p vs dc11.eff_p dc12.id_w_p vs dc12.eff_p dc13.id_w_p vs dc13.eff_p dc14.id_w_p vs dc14.eff_p

plot dc1.eff_ft_p vs dc1.eff_p dc2.eff_ft_p vs dc2.eff_p dc3.eff_ft_p vs dc3.eff_p dc4.eff_ft_p vs dc4.eff_p dc5.eff_ft_p vs dc5.eff_p dc6.eff_ft_p vs dc6.eff_p dc7.eff_ft_p vs dc7.eff_p dc8.eff_ft_p vs dc8.eff_p dc9.eff_ft_p vs dc9.eff_p dc10.eff_ft_p vs dc10.eff_p dc11.eff_ft_p vs dc11.eff_p dc12.eff_ft_p vs dc12.eff_p dc13.eff_ft_p vs dc13.eff_p dc14.eff_ft_p vs dc14.eff_p
.endc
